module block_gen # (
    parameter Param0,
    parameter Param1,
    parameter Param2
)  (
    input logic Port0,
    input logic Port1,
    input logic Port2
);

endmodule: block_gen

