interface test_if_params_array # (
    parameter param1,
    parameter param2
)   (
    input logic clk,
    input logic rst_n
);

endinterface: test_if_params_array

