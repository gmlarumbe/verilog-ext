`ifndef <UVM_NAME>_TYPES
`define <UVM_NAME>_TYPES

typedef enum bit {FALSE=0, TRUE=1} bool_t;

`endif // <UVM_NAME>_TYPES
