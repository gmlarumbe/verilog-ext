module foo # (
parameter integer A = 0,
B = 0,
C = 10,
parameter D = 0,
F = 0,
parameter int G = 0,
H = 1,
J = 0
)(
input wire a,
input wire b,
output reg z
);
endmodule


// Local Variables:
// verilog-indent-lists: nil
// End:
