
module x;

    foo;
endmodule

bar;
module z;
endmodule
