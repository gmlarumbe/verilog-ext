module foo
// ...
function asdf;
    // ...
endfunction
// ...
task asdf;
    // ...
endtask
// ...
generate
    // ...
    endgenerate
    // ...
covergroup
    // ...
    endgroup
    // ...
    property
    // ...
endproperty
// ...
sequence
    // ...
    endsequence
    // ...
    endmodule
// ...

// ...
package foo;
    // ...
    class foo2;
        // ...
    endclass
    // ...
endpackage
// ...

class foo3;
    // ...
endclass
// ...

virtual class foo4;
    // ...
endclass
// ...

interface class foo5;
    // ...
endclass
// ...

class foo6;
    // ...
    class foo7;
        // ...
    endclass
    // ...
endclass
// ...

program
    // ...
    endprogram
// ...
