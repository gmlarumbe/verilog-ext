`ifndef <UVM_NAME>_TYPES
`define <UVM_NAME>_TYPES



`endif // <UVM_NAME>_TYPES
