module block1 (
    input logic Port0,
    input logic Port1,
    input logic Port2
);

endmodule: block1

