module foo(reg_input_signal_name);
    input a;
    input    reg_input_signal_name;

endmodule // foo

