
module x;

    foo foo;
endmodule

bar bar;
module z;
endmodule
