interface test_if_params_empty (
    input logic clk,
    input logic rst_n
);

endinterface: test_if_params_empty

