interface <uvm_name>_if #(
    // ...
) ();

    logic clk;
    logic resetn;

    // ...

endinterface

