interface test_if (
    input logic clk,
    input logic rst_n
);

endinterface: test_if

